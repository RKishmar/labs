library verilog;
use verilog.vl_types.all;
entity lab2_6_tb is
end lab2_6_tb;
