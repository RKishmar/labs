
logic [$clog2($data_i(N)+1)-1:0] data_o;
